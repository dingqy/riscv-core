module RegisterFile(
  
);



endmodule // 