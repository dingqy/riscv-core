module Digit(
  input [31:0] data,
  input AN
);

endmodule // 